//=========================================================================
// Name & Email must be EXACTLY as in Gradescope roster!
// Name: Nicole Navarro 
// Email: nnava026@ucr.edu
// 
// Assignment name: Lab 3 Carry Look Ahead Adder
// Lab section: 021
// TA: Jincong Lu
// 
// I hereby certify that I have not received assistance on this assignment,
// or used code, from ANY outside source other than the instruction team
// (apart from what was provided in the starter file).
//
//=========================================================================

`timescale 1ns / 1ps

//  Constant definitions 

module carry_look_ahead_adder # ( parameter NUMBITS = 16 ) (
  input  wire[NUMBITS-1:0] A, 
  input  wire[NUMBITS-1:0] B, 
  input wire carryin, 
  output reg [NUMBITS-1:0] result,  
  output reg carryout
);

    // ------------------------------
    // Insert your solution below
    // ------------------------------ 

endmodule